//0616087
//Subject:     CO project 4 - Adder
//--------------------------------------------------------------------------------
//Version:     1
//--------------------------------------------------------------------------------
//Writer:      perry
//----------------------------------------------
//Date:        
//----------------------------------------------
//Description: 
//--------------------------------------------------------------------------------

module Adder(
    src1_i,
	src2_i,
	sum_o
	);

input  [32-1:0]  src1_i;
input  [32-1:0]	 src2_i;
output [32-1:0]	 sum_o;

wire   [32-1:0]	 sum_o;

reg    [32-1:0]  result;

always@(*)begin
    result = {src1_i + src2_i};
end

assign sum_o = result;

endmodule